// Verilog test fixture created from schematic C:\Users\Elizabeth\Documents\CE 1202 Lab\ToyProcessor\nor8.sch - Wed Jan 25 16:35:51 2017

`timescale 1ns / 1ps

module nor8_nor8_sch_tb();

// Inputs
   reg [7:0] zero_in;

// Output
   wire zero_out;

// Bidirs


endmodule
