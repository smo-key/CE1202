// Verilog Test Fixture Template

`timescale 1 ns / 1 ps

module mux_2to1_8bit_vtest();
	
endmodule
